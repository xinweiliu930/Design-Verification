module module4SVA (
input clk, quick_n_reset, i_wb_ack, extra_write_r,[2:0] wishbone_st
);

import FSMProperties::*;

// states recreated
localparam [3:0] WB_IDLE            = 3'd0,
                 WB_BURST1          = 3'd1,
                 WB_BURST2          = 3'd2,
                 WB_BURST3          = 3'd3,
                 WB_WAIT_ACK        = 3'd4;


/*place your properties here*/

assert property(FSMValidTransition(wishbone_st == WB_IDLE,1, wishbone_st == WB_IDLE||wishbone_st == WB_BURST1 || wishbone_st == WB_WAIT_ACK,clk,quick_n_reset ));
assert property(FSMValidTransition(wishbone_st == WB_BURST1,i_wb_ack, wishbone_st == WB_BURST2,clk,quick_n_reset));
assert property(FSMValidTransition(wishbone_st == WB_BURST2,i_wb_ack,wishbone_st == WB_BURST3 ,clk,quick_n_reset));
assert property(FSMValidTransition(wishbone_st == WB_BURST3,i_wb_ack,wishbone_st == WB_WAIT_ACK ,clk,quick_n_reset));
assert property(FSMValidTransition(wishbone_st == WB_WAIT_ACK,extra_write_r||!i_wb_ack, wishbone_st == WB_WAIT_ACK,clk,quick_n_reset));
assert property(FSMValidTransition(wishbone_st == WB_WAIT_ACK,!extra_write_r&&i_wb_ack,wishbone_st == WB_IDLE,clk,quick_n_reset));
assert property(FSMTimeOut(wishbone_st,1000,clk,quick_n_reset));


endmodule

module Wrapper ;

bind a25_wishbone module4SVA wrp (

.clk(i_clk),
.quick_n_reset(quick_n_reset),
.i_wb_ack(i_wb_ack),
.extra_write_r(extra_write_r),
.wishbone_st(wishbone_st));

endmodule
